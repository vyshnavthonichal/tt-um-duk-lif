magic
tech sky130A
magscale 1 2
timestamp 1713507025
<< locali >>
rect 22141 8637 22235 8642
rect 22141 8558 22239 8637
rect 22141 8381 22235 8558
rect 22141 8324 22157 8381
rect 22220 8324 22235 8381
rect 22141 8305 22235 8324
<< viali >>
rect 22157 8324 22220 8381
<< metal1 >>
rect 2256 12118 2706 12196
rect 2256 12096 25346 12118
rect 2256 11820 2340 12096
rect 2636 11820 25346 12096
rect 2256 11813 25346 11820
rect 2256 11704 2706 11813
rect 25041 9453 25346 11813
rect 26063 8790 26692 8808
rect 26063 8779 26594 8790
rect 26574 8698 26594 8779
rect 26676 8698 26692 8790
rect 26574 8678 26692 8698
rect 22141 8381 22235 8400
rect 22141 8324 22157 8381
rect 22220 8324 22235 8381
rect 22141 8305 22235 8324
rect 26276 8016 26408 8040
rect 26276 7930 26304 8016
rect 25903 7922 26304 7930
rect 26388 7922 26408 8016
rect 25903 7889 26408 7922
rect 26276 7888 26408 7889
rect 11360 5127 11710 5206
rect 24469 5127 24759 7377
rect 11360 5114 24759 5127
rect 11360 4876 11414 5114
rect 11656 4876 24759 5114
rect 11360 4837 24759 4876
rect 11360 4778 11710 4837
<< via1 >>
rect 2340 11820 2636 12096
rect 26594 8698 26676 8790
rect 26304 7922 26388 8016
rect 11414 4876 11656 5114
<< metal2 >>
rect 2256 12096 2706 12196
rect 2256 11820 2340 12096
rect 2636 11820 2706 12096
rect 2256 11704 2706 11820
rect 26574 8790 26692 8808
rect 26574 8698 26594 8790
rect 26676 8698 26692 8790
rect 26574 8678 26692 8698
rect 22141 8305 22235 8400
rect 11360 5114 11710 5206
rect 11360 4876 11414 5114
rect 11656 4876 11710 5114
rect 11360 4778 11710 4876
rect 22157 4512 22220 8305
rect 26276 8016 26408 8040
rect 26276 7922 26304 8016
rect 26388 7922 26408 8016
rect 26276 7888 26408 7922
rect 22136 4407 22646 4512
rect 22541 3895 22646 4407
rect 22480 3860 22647 3895
rect 22480 3695 22500 3860
rect 22626 3695 22647 3860
rect 22480 3666 22647 3695
<< via2 >>
rect 2340 11820 2636 12096
rect 26594 8698 26676 8790
rect 11414 4876 11656 5114
rect 26304 7922 26388 8016
rect 22500 3695 22626 3860
<< metal3 >>
rect 2256 12096 2706 12196
rect 2256 11820 2340 12096
rect 2636 11820 2706 12096
rect 2256 11704 2706 11820
rect 26574 8790 26692 8808
rect 26574 8698 26594 8790
rect 26676 8698 26692 8790
rect 26574 8678 26692 8698
rect 26276 8016 26408 8040
rect 26276 7922 26304 8016
rect 26388 7922 26408 8016
rect 26276 7888 26408 7922
rect 11360 5114 11710 5206
rect 11360 4876 11414 5114
rect 11656 4876 11710 5114
rect 11360 4778 11710 4876
rect 22480 3860 22647 3895
rect 22480 3695 22500 3860
rect 22626 3695 22647 3860
rect 22480 3666 22647 3695
<< via3 >>
rect 2340 11820 2636 12096
rect 26594 8698 26676 8790
rect 26304 7922 26388 8016
rect 11414 4876 11656 5114
rect 22500 3695 22626 3860
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 12080 500 44152
rect 2256 12096 2706 12196
rect 2256 12080 2340 12096
rect 200 11820 2340 12080
rect 2636 11820 2706 12096
rect 200 11808 2706 11820
rect 200 1000 500 11808
rect 2256 11704 2706 11808
rect 9800 5092 10100 44152
rect 26574 8798 26692 8808
rect 26574 8790 31432 8798
rect 26574 8698 26594 8790
rect 26676 8698 31432 8790
rect 26574 8678 31432 8698
rect 26276 8016 27016 8040
rect 26276 7922 26304 8016
rect 26388 7922 27016 8016
rect 26276 7920 27016 7922
rect 26276 7888 26408 7920
rect 11360 5114 11710 5206
rect 11360 5092 11414 5114
rect 9800 4876 11414 5092
rect 11656 4876 11710 5114
rect 9800 4868 11710 4876
rect 9800 1000 10100 4868
rect 11360 4778 11710 4868
rect 22480 3860 22647 3895
rect 22480 3695 22500 3860
rect 22626 3695 22647 3860
rect 22480 3666 22647 3695
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 3666
rect 26896 0 27016 7920
rect 31312 0 31432 8678
use leakylayout  leakylayout_0 ~/Desktop/tt_vyshnav/new/leaky.sch
timestamp 1713507025
transform 1 0 22750 0 1 6922
box -6156 -3517 3342 3488
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
