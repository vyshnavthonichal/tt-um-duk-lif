VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_duk_lif
  CLASS BLOCK ;
  FOREIGN tt_um_duk_lif ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.976400 ;
    ANTENNADIFFAREA 28.198374 ;
    PORT
      LAYER nwell ;
        RECT 110.800 44.260 126.530 47.210 ;
        RECT 114.370 44.075 115.245 44.260 ;
        RECT 119.155 44.055 126.530 44.260 ;
        RECT 119.155 42.525 126.515 44.055 ;
        RECT 119.155 42.045 126.510 42.525 ;
        RECT 119.155 41.850 126.490 42.045 ;
        RECT 119.155 41.820 124.860 41.850 ;
        RECT 123.365 41.785 124.860 41.820 ;
        RECT 123.365 41.760 124.795 41.785 ;
      LAYER li1 ;
        RECT 111.105 45.190 114.355 48.660 ;
        RECT 115.330 45.195 118.580 48.660 ;
        RECT 111.090 45.020 114.370 45.190 ;
        RECT 115.320 45.025 118.600 45.195 ;
        RECT 119.790 45.190 123.040 48.660 ;
        RECT 115.320 44.555 118.600 44.725 ;
        RECT 119.175 44.650 119.510 45.075 ;
        RECT 119.770 45.020 123.050 45.190 ;
        RECT 124.410 45.185 125.610 48.660 ;
        RECT 124.390 45.015 125.630 45.185 ;
        RECT 116.495 43.950 116.875 44.555 ;
        RECT 116.495 43.935 118.695 43.950 ;
        RECT 116.495 43.700 118.705 43.935 ;
        RECT 118.490 42.930 118.705 43.700 ;
        RECT 115.190 42.355 115.650 42.835 ;
        RECT 115.870 42.760 118.710 42.930 ;
        RECT 118.490 41.605 118.705 42.760 ;
        RECT 119.275 42.565 119.445 44.650 ;
        RECT 119.770 44.550 123.050 44.720 ;
        RECT 120.135 44.270 122.930 44.550 ;
        RECT 124.390 44.545 125.630 44.715 ;
        RECT 124.885 44.350 125.055 44.545 ;
        RECT 120.135 44.100 124.005 44.270 ;
        RECT 124.880 44.145 125.055 44.350 ;
        RECT 120.135 43.910 122.930 44.100 ;
        RECT 119.880 42.700 123.120 43.910 ;
        RECT 123.835 43.515 124.005 44.100 ;
        RECT 124.815 43.805 125.140 44.145 ;
        RECT 123.835 43.510 125.345 43.515 ;
        RECT 123.835 43.345 125.355 43.510 ;
        RECT 124.555 42.920 125.355 43.345 ;
        RECT 127.445 43.215 127.890 43.585 ;
        RECT 127.550 42.980 127.760 43.215 ;
        RECT 124.535 42.750 125.375 42.920 ;
        RECT 126.985 42.810 128.525 42.980 ;
        RECT 119.180 42.170 119.555 42.565 ;
        RECT 119.860 42.530 123.140 42.700 ;
        RECT 119.290 41.605 119.460 42.170 ;
        RECT 118.490 41.425 119.465 41.605 ;
        RECT 118.505 41.420 119.465 41.425 ;
        RECT 119.290 41.175 119.460 41.420 ;
        RECT 120.085 41.175 120.390 41.255 ;
        RECT 119.290 41.150 120.390 41.175 ;
        RECT 119.285 41.005 120.390 41.150 ;
        RECT 119.285 38.795 119.460 41.005 ;
        RECT 120.085 40.900 120.390 41.005 ;
        RECT 120.205 38.795 120.545 38.890 ;
        RECT 119.285 38.620 120.545 38.795 ;
        RECT 119.285 34.755 119.500 38.620 ;
        RECT 120.205 38.540 120.545 38.620 ;
        RECT 118.465 33.585 120.130 34.755 ;
        RECT 85.405 30.105 88.605 30.860 ;
        RECT 85.405 28.695 92.135 30.105 ;
        RECT 85.405 28.070 88.605 28.695 ;
      LAYER mcon ;
        RECT 112.305 47.580 113.140 48.335 ;
        RECT 116.580 47.570 117.415 48.325 ;
        RECT 120.970 47.565 121.805 48.320 ;
        RECT 111.170 45.020 114.290 45.190 ;
        RECT 115.400 45.025 118.520 45.195 ;
        RECT 124.615 47.545 125.450 48.300 ;
        RECT 115.400 44.555 118.520 44.725 ;
        RECT 119.850 45.020 122.970 45.190 ;
        RECT 124.470 45.015 125.550 45.185 ;
        RECT 115.250 42.440 115.600 42.770 ;
        RECT 115.950 42.760 117.330 42.930 ;
        RECT 119.850 44.550 122.970 44.720 ;
        RECT 124.470 44.545 125.550 44.715 ;
        RECT 124.875 43.860 125.075 44.070 ;
        RECT 127.575 43.305 127.785 43.490 ;
        RECT 124.615 42.750 125.295 42.920 ;
        RECT 127.065 42.810 128.445 42.980 ;
        RECT 119.940 42.530 123.060 42.700 ;
        RECT 118.780 33.735 119.795 34.570 ;
        RECT 86.220 28.720 87.980 30.215 ;
        RECT 90.065 28.775 92.050 30.025 ;
      LAYER met1 ;
        RECT 11.280 60.590 13.530 60.980 ;
        RECT 11.280 59.065 126.730 60.590 ;
        RECT 11.280 58.520 13.530 59.065 ;
        RECT 125.205 48.660 126.730 59.065 ;
        RECT 110.800 47.265 126.730 48.660 ;
        RECT 110.800 47.260 126.485 47.265 ;
        RECT 115.325 46.530 129.175 46.715 ;
        RECT 115.330 45.675 115.495 46.530 ;
        RECT 115.335 45.225 115.495 45.675 ;
        RECT 111.110 44.990 114.350 45.220 ;
        RECT 115.335 44.995 118.580 45.225 ;
        RECT 115.335 44.755 115.495 44.995 ;
        RECT 119.790 44.990 123.030 45.220 ;
        RECT 124.410 44.985 125.610 45.215 ;
        RECT 115.335 44.525 118.580 44.755 ;
        RECT 115.335 42.920 115.495 44.525 ;
        RECT 119.790 44.520 123.030 44.750 ;
        RECT 124.410 44.515 125.610 44.745 ;
        RECT 124.815 44.040 125.140 44.145 ;
        RECT 129.005 44.040 129.175 46.530 ;
        RECT 124.815 43.900 133.460 44.040 ;
        RECT 124.815 43.895 129.175 43.900 ;
        RECT 129.525 43.895 133.460 43.900 ;
        RECT 124.815 43.805 125.140 43.895 ;
        RECT 127.600 43.585 127.740 43.895 ;
        RECT 127.445 43.215 127.890 43.585 ;
        RECT 132.870 43.390 133.460 43.895 ;
        RECT 115.110 42.255 115.725 42.920 ;
        RECT 115.890 42.730 117.390 42.960 ;
        RECT 119.880 42.500 123.120 42.730 ;
        RECT 124.555 42.720 125.355 42.950 ;
        RECT 127.005 42.780 128.505 43.010 ;
        RECT 115.335 42.250 115.550 42.255 ;
        RECT 118.465 33.585 120.130 34.755 ;
        RECT 85.405 28.070 88.605 30.860 ;
        RECT 90.005 28.745 92.110 30.055 ;
      LAYER via ;
        RECT 11.700 59.100 13.180 60.480 ;
        RECT 132.970 43.490 133.380 43.950 ;
        RECT 118.780 33.735 119.795 34.570 ;
        RECT 86.220 28.720 87.980 30.215 ;
      LAYER met2 ;
        RECT 11.280 58.520 13.530 60.980 ;
        RECT 132.870 43.390 133.460 44.040 ;
        RECT 118.465 33.585 120.130 34.755 ;
        RECT 85.405 28.070 88.605 30.860 ;
      LAYER via2 ;
        RECT 11.700 59.100 13.180 60.480 ;
        RECT 132.970 43.490 133.380 43.950 ;
        RECT 118.780 33.735 119.795 34.570 ;
        RECT 86.220 28.720 87.980 30.215 ;
      LAYER met3 ;
        RECT 11.280 58.520 13.530 60.980 ;
        RECT 132.870 43.390 133.460 44.040 ;
        RECT 118.465 33.585 120.130 34.755 ;
        RECT 85.405 28.070 88.605 30.860 ;
      LAYER via3 ;
        RECT 11.700 59.100 13.180 60.480 ;
        RECT 132.970 43.490 133.380 43.950 ;
        RECT 118.780 33.735 119.795 34.570 ;
        RECT 86.220 28.720 87.980 30.215 ;
      LAYER met4 ;
        RECT 1.000 60.400 2.500 220.760 ;
        RECT 11.280 60.400 13.530 60.980 ;
        RECT 1.000 59.040 13.530 60.400 ;
        RECT 1.000 5.000 2.500 59.040 ;
        RECT 11.280 58.520 13.530 59.040 ;
        RECT 83.365 32.045 107.975 51.655 ;
        RECT 132.870 43.990 133.460 44.040 ;
        RECT 132.870 43.390 157.160 43.990 ;
        RECT 118.465 33.585 120.130 34.755 ;
        RECT 86.200 30.860 87.615 32.045 ;
        RECT 107.015 31.145 107.975 32.045 ;
        RECT 118.780 31.145 119.800 33.585 ;
        RECT 107.015 31.130 119.800 31.145 ;
        RECT 85.405 28.070 88.605 30.860 ;
        RECT 107.015 30.330 119.765 31.130 ;
        RECT 156.560 0.000 157.160 43.390 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 125.080 39.335 125.525 39.705 ;
        RECT 125.185 39.040 125.405 39.335 ;
        RECT 124.540 38.870 126.080 39.040 ;
      LAYER mcon ;
        RECT 125.195 39.415 125.390 39.640 ;
        RECT 124.620 38.870 126.000 39.040 ;
      LAYER met1 ;
        RECT 125.080 39.650 125.525 39.705 ;
        RECT 131.380 39.650 132.040 40.200 ;
        RECT 125.080 39.445 132.040 39.650 ;
        RECT 125.080 39.335 125.525 39.445 ;
        RECT 131.380 39.440 132.040 39.445 ;
        RECT 124.560 38.840 126.060 39.070 ;
      LAYER via ;
        RECT 131.520 39.610 131.940 40.080 ;
      LAYER met2 ;
        RECT 131.380 39.440 132.040 40.200 ;
      LAYER via2 ;
        RECT 131.520 39.610 131.940 40.080 ;
      LAYER met3 ;
        RECT 131.380 39.440 132.040 40.200 ;
      LAYER via3 ;
        RECT 131.520 39.610 131.940 40.080 ;
      LAYER met4 ;
        RECT 131.380 39.600 135.080 40.200 ;
        RECT 131.380 39.440 132.040 39.600 ;
        RECT 134.480 0.000 135.080 39.600 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.705 41.525 111.175 42.000 ;
        RECT 110.785 22.560 111.100 41.525 ;
        RECT 110.680 22.035 113.230 22.560 ;
        RECT 112.705 19.475 113.230 22.035 ;
        RECT 112.400 18.330 113.235 19.475 ;
      LAYER via2 ;
        RECT 112.500 18.475 113.130 19.300 ;
      LAYER met3 ;
        RECT 112.400 18.330 113.235 19.475 ;
      LAYER via3 ;
        RECT 112.500 18.475 113.130 19.300 ;
      LAYER met4 ;
        RECT 112.400 18.330 113.235 19.475 ;
        RECT 112.400 0.000 113.000 18.330 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 111.720 42.665 113.760 42.835 ;
        RECT 111.740 41.930 113.740 42.665 ;
        RECT 115.870 42.290 117.410 42.460 ;
        RECT 111.750 36.320 113.740 41.930 ;
        RECT 115.885 41.330 117.390 42.290 ;
        RECT 124.535 42.280 125.375 42.450 ;
        RECT 126.985 42.340 128.525 42.510 ;
        RECT 124.870 41.625 125.040 42.280 ;
        RECT 115.940 36.320 117.300 41.330 ;
        RECT 124.800 41.275 125.145 41.625 ;
        RECT 127.005 41.510 128.505 42.340 ;
        RECT 120.760 38.385 122.300 38.555 ;
        RECT 120.780 37.560 122.280 38.385 ;
        RECT 120.790 36.320 122.275 37.560 ;
        RECT 127.010 36.320 128.500 41.510 ;
        RECT 115.430 33.565 117.220 34.715 ;
        RECT 115.635 33.315 117.050 33.565 ;
        RECT 115.630 32.280 117.050 33.315 ;
        RECT 111.155 30.865 129.495 32.280 ;
        RECT 128.080 30.105 129.495 30.865 ;
        RECT 127.575 28.695 129.735 30.105 ;
      LAYER mcon ;
        RECT 111.800 42.665 113.680 42.835 ;
        RECT 115.950 42.290 117.330 42.460 ;
        RECT 124.615 42.280 125.295 42.450 ;
        RECT 127.065 42.340 128.445 42.510 ;
        RECT 124.880 41.350 125.055 41.525 ;
        RECT 112.045 36.510 113.410 36.915 ;
        RECT 120.840 38.385 122.220 38.555 ;
        RECT 116.240 36.560 117.010 36.950 ;
        RECT 120.945 36.510 122.095 36.930 ;
        RECT 127.435 36.525 128.135 36.980 ;
        RECT 115.780 33.760 116.885 34.535 ;
        RECT 127.660 28.775 129.645 30.025 ;
      LAYER met1 ;
        RECT 111.740 42.635 113.740 42.865 ;
        RECT 115.890 42.260 117.390 42.490 ;
        RECT 124.555 42.250 125.355 42.480 ;
        RECT 127.005 42.310 128.505 42.540 ;
        RECT 124.800 41.275 125.145 41.625 ;
        RECT 124.855 41.090 125.095 41.275 ;
        RECT 123.590 40.850 125.095 41.090 ;
        RECT 120.780 38.355 122.280 38.585 ;
        RECT 123.590 37.100 123.830 40.850 ;
        RECT 110.950 36.320 128.510 37.100 ;
        RECT 115.835 34.940 116.885 36.320 ;
        RECT 115.430 33.565 117.220 34.940 ;
        RECT 56.800 25.635 58.550 26.030 ;
        RECT 122.345 25.635 123.795 36.320 ;
        RECT 127.600 28.745 129.705 30.055 ;
        RECT 56.800 24.185 123.795 25.635 ;
        RECT 56.800 23.890 58.550 24.185 ;
      LAYER via ;
        RECT 115.780 33.760 116.885 34.535 ;
        RECT 57.070 24.380 58.280 25.570 ;
      LAYER met2 ;
        RECT 115.430 33.565 117.220 34.715 ;
        RECT 56.800 23.890 58.550 26.030 ;
      LAYER via2 ;
        RECT 115.780 33.760 116.885 34.535 ;
        RECT 57.070 24.380 58.280 25.570 ;
      LAYER met3 ;
        RECT 82.970 34.275 109.830 52.050 ;
        RECT 115.430 34.275 117.220 34.715 ;
        RECT 82.970 33.860 117.220 34.275 ;
        RECT 82.970 31.650 109.830 33.860 ;
        RECT 115.430 33.565 117.220 33.860 ;
        RECT 56.800 23.890 58.550 26.030 ;
      LAYER via3 ;
        RECT 109.410 31.790 109.730 51.910 ;
        RECT 57.070 24.380 58.280 25.570 ;
      LAYER met4 ;
        RECT 49.000 25.460 50.500 220.760 ;
        RECT 109.330 31.710 109.810 51.990 ;
        RECT 56.800 25.460 58.550 26.030 ;
        RECT 49.000 24.340 58.550 25.460 ;
        RECT 49.000 5.000 50.500 24.340 ;
        RECT 56.800 23.890 58.550 24.340 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 125.945 44.985 126.275 45.050 ;
        RECT 126.570 44.985 126.780 44.990 ;
        RECT 125.945 44.815 126.780 44.985 ;
        RECT 111.090 44.550 114.370 44.720 ;
        RECT 125.945 44.710 126.275 44.815 ;
        RECT 111.805 43.955 113.685 44.550 ;
        RECT 114.650 44.140 114.985 44.415 ;
        RECT 114.710 43.955 114.925 44.140 ;
        RECT 111.805 43.770 114.925 43.955 ;
        RECT 111.805 43.305 113.685 43.770 ;
        RECT 126.570 43.420 126.780 44.815 ;
        RECT 110.705 43.185 111.175 43.210 ;
        RECT 110.705 42.790 111.495 43.185 ;
        RECT 111.720 43.135 113.760 43.305 ;
        RECT 125.900 43.250 126.780 43.420 ;
        RECT 110.705 41.525 111.175 42.790 ;
        RECT 124.045 42.430 124.360 42.765 ;
        RECT 119.860 42.060 123.140 42.230 ;
        RECT 120.760 41.780 122.140 42.060 ;
        RECT 120.760 41.605 122.965 41.780 ;
        RECT 120.760 41.405 122.140 41.605 ;
        RECT 120.710 41.235 122.250 41.405 ;
        RECT 122.795 41.240 122.965 41.605 ;
        RECT 122.795 41.050 122.970 41.240 ;
        RECT 120.710 40.765 122.250 40.935 ;
        RECT 120.730 39.960 122.230 40.765 ;
        RECT 122.800 40.680 122.970 41.050 ;
        RECT 124.115 40.680 124.295 42.430 ;
        RECT 125.900 40.680 126.130 43.250 ;
        RECT 126.570 42.880 126.780 43.250 ;
        RECT 126.430 42.480 126.800 42.880 ;
        RECT 122.800 40.510 126.130 40.680 ;
        RECT 120.875 39.595 122.090 39.960 ;
        RECT 120.875 39.585 123.495 39.595 ;
        RECT 120.875 39.415 123.500 39.585 ;
        RECT 120.875 39.025 122.090 39.415 ;
        RECT 120.760 38.855 122.300 39.025 ;
        RECT 123.295 37.930 123.500 39.415 ;
        RECT 124.115 38.915 124.305 40.510 ;
        RECT 124.515 40.505 125.935 40.510 ;
        RECT 124.085 38.535 124.360 38.915 ;
        RECT 124.540 38.400 126.080 38.570 ;
        RECT 124.555 37.930 126.065 38.400 ;
        RECT 123.295 37.745 126.065 37.930 ;
        RECT 124.555 37.560 126.065 37.745 ;
      LAYER mcon ;
        RECT 111.170 44.550 114.290 44.720 ;
        RECT 111.800 43.135 113.680 43.305 ;
        RECT 119.940 42.060 123.060 42.230 ;
        RECT 110.785 41.620 111.100 41.905 ;
        RECT 120.790 41.235 122.170 41.405 ;
        RECT 120.790 40.765 122.170 40.935 ;
        RECT 120.840 38.855 122.220 39.025 ;
        RECT 124.620 38.400 126.000 38.570 ;
      LAYER met1 ;
        RECT 111.110 44.520 114.350 44.750 ;
        RECT 111.740 43.105 113.740 43.335 ;
        RECT 119.880 42.030 123.120 42.260 ;
        RECT 110.705 41.525 111.175 42.000 ;
        RECT 120.730 41.205 122.230 41.435 ;
        RECT 120.730 40.735 122.230 40.965 ;
        RECT 120.780 38.825 122.280 39.055 ;
        RECT 124.560 38.370 126.060 38.600 ;
  END
END tt_um_duk_lif
END LIBRARY

